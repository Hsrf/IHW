module ControlUnit(
	input clock,
	input wire opcode [5:0],
	output wire pcWriteCond [1:0],
	output wire pcWrite [1:0],
	output wire iord [3:0],
	output wire memRead [1:0],
	output wire memWrite [1:0],
	output wire irWrite [1:0],
	output wire regDst [2:0],
	output wire regWrite [1:0],
	output wire writeRegA [1:0],
	output wire writeRegB [1:0],
	output wire aluSrcA [2:0],
	output wire aluSrcB [3:0],
	output wire aluOutControl [1:0],
	output wire epcWrite [1:0],
	output wire pcSource [3:0],
	output wire memToReg [4:0],
	output wire aluOp [3:0],
	output wire sControl [2:0],
	output wire memMux [1:0],
	output wire lsControl [2:0],
	output wire multControl [1:0],
	output wire divControl [1:0],
	output wire muxHiControl [1:0],
	output wire muxLoControl [1:0],
	output wire writeHI [1:0],
	output wire writeLO [1:0],
	output wire shiftSrc [1:0],
	output wire shiftAmt [1:0],
	output wire shiftControl [3:0],
	output wire divZero [1:0],
	output wire overflow [1:0]
);